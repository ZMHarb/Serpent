library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use work.mypackage.all;

entity tb_key_schedule is
end entity tb_key_schedule;

architecture Behavioral of tb_key_schedule is

    signal key_in_tb    : std_logic_vector(255 downto 0);
    signal roundkeys_tb : array_33x128;
    
    signal cmp_roundkeys : array_33x128 := 
(
 "01101111110001000111100001101001110100110101001101011001001110001000110101110101101111011001000011011111110110101000100101100111",
 "00010101101100100010101100111011111001101001001011101110011010001011110111111010000101100010110010010100110110111011011010010111",
 "00101101011000011111011111010100111000101011000010000111010111101010100100011010111110000001010100010010001111001000010000011010",
 "10001010000000110011010010100001010110110001100000010100100110000111100110111111100001011000111110000011000110110110110001010001",
 "10010110101010111011100111011000001101000110011111001001110111111010101101101111000111100001010010100111100010000101011111010011",
 "10111010101001001100100011010111000110100011010010111101100101010101110001011010100111001011111110111101100011101110101010010101",
 "01010010000010011011100000010001011001000000010101100000100000100010001000101011010100010001111010001100111101000001110101101000",
 "10110101001011001010000111101100010000001110110101010111100010100100101000101101001101010010111110111011101100101100111010000110",
 "10000000011100111110100110011101011110110011110101000111011011001000110101100000010000101111100111101110100100111011110011010011",
 "00111000001000110000100111000110000101101100101000001110110011101100010010011010011111010001110101001011011010001100001101110100",
 "10001110010001101000011010100100001001110101000000001000100101100111111000010101001010000000110110010001011111010001111101100100",
 "11101110100011101010110010011011000001010111000001001001111101001110110100010110101110110010010101010110100010001100010111001010",
 "11001101001111110001000111110110100101011111101101001011001001110110111010010111011001001100011101000111110111001011011011011000",
 "10110111100000001110100111000000001111110000110010110111010001010011011110010111011110001010001100111110101101011100111100000000",
 "10100101011011001100001110101100010011000011101110111100111110000010010111011101010010110001111010100101000010111010000110001111",
 "10101010110111101011000000000111010000100101100001100000000011110110100100110100101001111001010111001001011111111101010011101010",
 "11101001001000111100110000110010000100000101111101011110100110000110101000110110101111101011110011101001011001001000101001000100",
 "00010111011000000101000111001010110101001111000110110110111000011111101111011001110110011101111111010101010101101011100110110001",
 "01100110100000010101010011001001100011110111001100111000000000110110101101010011100010011001101100111011010001100101111100010001",
 "01011110111111100010011100111011001100010001111111000011110111000010110111001100010100001011010100001000111110000000100100011001",
 "10000001001110000011101010111011111100110110111110011110001100000111111101000011010001100110010010100000011000110011011100011000",
 "01001011000000111010110101111100100101000001111101001111011000101000101011010101111101000110100010000001001010001010011010111000",
 "10001101100100010010001110010001001111110101101000001000000100100001001101101011110010010101111101000101110101011011100111001010",
 "11111000011110010111011010010111011000101101110111011001010001011100111111001001000010000101011000000101111101000101010101001000",
 "11101111000111010000010000010011010111100000001010011001101001101010101100001110110101000111001001010101010010100100001100000010",
 "01000001111101011010000100000100110000110010010010101110001001001111110101000100110010111101110110101110100100011000011101011111",
 "10111011000100110010111010100011101001011010111000101111010111100000001011011001010011001110101000101001111100101011101101101110",
 "11110011001101100011100101000111101000010100111111011110101010010100100010000111111101001111100101100101011010010110011101010010",
 "00111001011110100110110011010000110011001000111010000011001110000101110000010111110101110010100101110000001001000111111100101010",
 "10100100101111010101101010010011111011000110100111011010011010001011001100100001010101100011010110110010111100000010011011111011",
 "11101101001110100111010110100001010101001000010101100110000011111100010100111010010111001101111110100001111111110010001000101111",
 "00101100011111111001011001101110110110001101010000110111101101100111110011000101101000011011011111000010011101100101101001000001",
 "10111001011101001000001101000010111000011011010001000101101111110111101110101100010111110010111001101010110001011110000110011001"
);

begin

    uut: entity work.key_schedule
        port map (
            key_in      => key_in_tb,
            round_keys  => roundkeys_tb
        );

    stim_proc: process
    begin

        key_in_tb <= x"00000000000000000000000000000001432da46b89ac716907cb7dcfcbcc9566";
        wait for 10ns;
        assert roundkeys_tb = cmp_roundkeys report "KeySchedule Error";

    end process;

end architecture Behavioral;
